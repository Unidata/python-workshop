netcdf mslp {
dimensions:
	lat = 6 ;
	lon = 4 ;
	time = UNLIMITED ; // (2 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
	double time(time) ;
		time:units = "seconds since 2009-01-01" ;
	float pr(time, lat, lon) ;
		pr:standard_name = "air_pressure_at_sea_level" ;
		pr:units = "hPa" ;

// global attributes:
		:title = "example for workshop updated" ;
data:

 lat = 25, 30, 35, 40, 45, 50 ;

 lon = -125, -110, -95, -80 ;

 time = 7776000, 15552000 ;

 pr =
  900.5, 901, 902, 903,
  904, 905, 906, 907,
  908, 909, 910, 911,
  912, 913, 914, 915,
  916, 917, 918, 919,
  920, 921, 922, 923,
  972, 973, 974, 975,
  976, 977, 978, 979,
  980, 981, 982, 983,
  984, 985, 986, 987,
  988, 989, 990, 991,
  992, 993, 994, 995 ;
}
